module verilog_module
  (
    input CLK,
    input c_en,
    output last_signal  
  );

always @(posedge CLK) begin
  # Set registers
end

endmodule
